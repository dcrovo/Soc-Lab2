-- nios2_p3.vhd

-- Generated using ACDS version 21.1 850

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios2_p3 is
	port (
		clk_clk       : in  std_logic                    := '0';             --    clk.clk
		hex_0_export  : out std_logic_vector(6 downto 0);                    --  hex_0.export
		hex_1_export  : out std_logic_vector(6 downto 0);                    --  hex_1.export
		hex_2_export  : out std_logic_vector(6 downto 0);                    --  hex_2.export
		hex_3_export  : out std_logic_vector(6 downto 0);                    --  hex_3.export
		hex_4_export  : out std_logic_vector(6 downto 0);                    --  hex_4.export
		hex_5_export  : out std_logic_vector(6 downto 0);                    --  hex_5.export
		reset_reset_n : in  std_logic                    := '0';             --  reset.reset_n
		switch_export : in  std_logic_vector(6 downto 0) := (others => '0')  -- switch.export
	);
end entity nios2_p3;

architecture rtl of nios2_p3 is
	component nios2_p3_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios2_p3_cpu;

	component nios2_p3_hex_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component nios2_p3_hex_0;

	component nios2_p3_onchip_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component nios2_p3_onchip_mem;

	component nios2_p3_switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(6 downto 0)  := (others => 'X')  -- export
		);
	end component nios2_p3_switch;

	component nios2_p3_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios2_p3_sysid;

	component nios2_p3_mm_interconnect_0 is
		port (
			clk_clk_clk                             : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			hex_5_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                 : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address          : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			hex_0_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_0_s1_write                          : out std_logic;                                        -- write
			hex_0_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_0_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_0_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_1_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_1_s1_write                          : out std_logic;                                        -- write
			hex_1_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_1_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_1_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_2_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_2_s1_write                          : out std_logic;                                        -- write
			hex_2_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_2_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_2_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_3_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_3_s1_write                          : out std_logic;                                        -- write
			hex_3_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_3_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_3_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_4_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_4_s1_write                          : out std_logic;                                        -- write
			hex_4_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_4_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_4_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_5_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_5_s1_write                          : out std_logic;                                        -- write
			hex_5_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_5_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_5_s1_chipselect                     : out std_logic;                                        -- chipselect
			onchip_mem_s1_address                   : out std_logic_vector(13 downto 0);                    -- address
			onchip_mem_s1_write                     : out std_logic;                                        -- write
			onchip_mem_s1_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem_s1_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem_s1_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem_s1_chipselect                : out std_logic;                                        -- chipselect
			onchip_mem_s1_clken                     : out std_logic;                                        -- clken
			switch_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			switch_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_control_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component nios2_p3_mm_interconnect_0;

	component nios2_p3_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios2_p3_irq_mapper;

	component nios2_p3_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios2_p3_rst_controller;

	component nios2_p3_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios2_p3_rst_controller_001;

	signal cpu_data_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                       : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                           : std_logic_vector(17 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                        : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                              : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                             : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                         : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                    : std_logic_vector(17 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                       : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_sysid_control_slave_readdata    : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata    : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read        : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write       : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_mem_s1_chipselect        : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	signal mm_interconnect_0_onchip_mem_s1_readdata          : std_logic_vector(31 downto 0); -- onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	signal mm_interconnect_0_onchip_mem_s1_address           : std_logic_vector(13 downto 0); -- mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	signal mm_interconnect_0_onchip_mem_s1_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	signal mm_interconnect_0_onchip_mem_s1_write             : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	signal mm_interconnect_0_onchip_mem_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	signal mm_interconnect_0_onchip_mem_s1_clken             : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	signal mm_interconnect_0_switch_s1_readdata              : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_s1_readdata
	signal mm_interconnect_0_switch_s1_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_s1_address -> switch:address
	signal mm_interconnect_0_hex_0_s1_chipselect             : std_logic;                     -- mm_interconnect_0:hex_0_s1_chipselect -> hex_0:chipselect
	signal mm_interconnect_0_hex_0_s1_readdata               : std_logic_vector(31 downto 0); -- hex_0:readdata -> mm_interconnect_0:hex_0_s1_readdata
	signal mm_interconnect_0_hex_0_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_0_s1_address -> hex_0:address
	signal mm_interconnect_0_hex_0_s1_write                  : std_logic;                     -- mm_interconnect_0:hex_0_s1_write -> mm_interconnect_0_hex_0_s1_write:in
	signal mm_interconnect_0_hex_0_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_0_s1_writedata -> hex_0:writedata
	signal mm_interconnect_0_hex_1_s1_chipselect             : std_logic;                     -- mm_interconnect_0:hex_1_s1_chipselect -> hex_1:chipselect
	signal mm_interconnect_0_hex_1_s1_readdata               : std_logic_vector(31 downto 0); -- hex_1:readdata -> mm_interconnect_0:hex_1_s1_readdata
	signal mm_interconnect_0_hex_1_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_1_s1_address -> hex_1:address
	signal mm_interconnect_0_hex_1_s1_write                  : std_logic;                     -- mm_interconnect_0:hex_1_s1_write -> mm_interconnect_0_hex_1_s1_write:in
	signal mm_interconnect_0_hex_1_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_1_s1_writedata -> hex_1:writedata
	signal mm_interconnect_0_hex_2_s1_chipselect             : std_logic;                     -- mm_interconnect_0:hex_2_s1_chipselect -> hex_2:chipselect
	signal mm_interconnect_0_hex_2_s1_readdata               : std_logic_vector(31 downto 0); -- hex_2:readdata -> mm_interconnect_0:hex_2_s1_readdata
	signal mm_interconnect_0_hex_2_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_2_s1_address -> hex_2:address
	signal mm_interconnect_0_hex_2_s1_write                  : std_logic;                     -- mm_interconnect_0:hex_2_s1_write -> mm_interconnect_0_hex_2_s1_write:in
	signal mm_interconnect_0_hex_2_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_2_s1_writedata -> hex_2:writedata
	signal mm_interconnect_0_hex_3_s1_chipselect             : std_logic;                     -- mm_interconnect_0:hex_3_s1_chipselect -> hex_3:chipselect
	signal mm_interconnect_0_hex_3_s1_readdata               : std_logic_vector(31 downto 0); -- hex_3:readdata -> mm_interconnect_0:hex_3_s1_readdata
	signal mm_interconnect_0_hex_3_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_3_s1_address -> hex_3:address
	signal mm_interconnect_0_hex_3_s1_write                  : std_logic;                     -- mm_interconnect_0:hex_3_s1_write -> mm_interconnect_0_hex_3_s1_write:in
	signal mm_interconnect_0_hex_3_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_3_s1_writedata -> hex_3:writedata
	signal mm_interconnect_0_hex_4_s1_chipselect             : std_logic;                     -- mm_interconnect_0:hex_4_s1_chipselect -> hex_4:chipselect
	signal mm_interconnect_0_hex_4_s1_readdata               : std_logic_vector(31 downto 0); -- hex_4:readdata -> mm_interconnect_0:hex_4_s1_readdata
	signal mm_interconnect_0_hex_4_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_4_s1_address -> hex_4:address
	signal mm_interconnect_0_hex_4_s1_write                  : std_logic;                     -- mm_interconnect_0:hex_4_s1_write -> mm_interconnect_0_hex_4_s1_write:in
	signal mm_interconnect_0_hex_4_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_4_s1_writedata -> hex_4:writedata
	signal mm_interconnect_0_hex_5_s1_chipselect             : std_logic;                     -- mm_interconnect_0:hex_5_s1_chipselect -> hex_5:chipselect
	signal mm_interconnect_0_hex_5_s1_readdata               : std_logic_vector(31 downto 0); -- hex_5:readdata -> mm_interconnect_0:hex_5_s1_readdata
	signal mm_interconnect_0_hex_5_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_5_s1_address -> hex_5:address
	signal mm_interconnect_0_hex_5_s1_write                  : std_logic;                     -- mm_interconnect_0:hex_5_s1_write -> mm_interconnect_0_hex_5_s1_write:in
	signal mm_interconnect_0_hex_5_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_5_s1_writedata -> hex_5:writedata
	signal cpu_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                    : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_mem:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                     : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:hex_5_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal reset_reset_n_ports_inv                           : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_hex_0_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_hex_0_s1_write:inv -> hex_0:write_n
	signal mm_interconnect_0_hex_1_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_hex_1_s1_write:inv -> hex_1:write_n
	signal mm_interconnect_0_hex_2_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_hex_2_s1_write:inv -> hex_2:write_n
	signal mm_interconnect_0_hex_3_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_hex_3_s1_write:inv -> hex_3:write_n
	signal mm_interconnect_0_hex_4_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_hex_4_s1_write:inv -> hex_4:write_n
	signal mm_interconnect_0_hex_5_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_hex_5_s1_write:inv -> hex_5:write_n
	signal rst_controller_reset_out_reset_ports_inv          : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, hex_0:reset_n, hex_1:reset_n, hex_2:reset_n, hex_3:reset_n, hex_4:reset_n, switch:reset_n, sysid:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv      : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> hex_5:reset_n

begin

	cpu : component nios2_p3_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	hex_0 : component nios2_p3_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_0_s1_readdata,        --                    .readdata
			out_port   => hex_0_export                                -- external_connection.export
		);

	hex_1 : component nios2_p3_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_1_s1_readdata,        --                    .readdata
			out_port   => hex_1_export                                -- external_connection.export
		);

	hex_2 : component nios2_p3_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_2_s1_readdata,        --                    .readdata
			out_port   => hex_2_export                                -- external_connection.export
		);

	hex_3 : component nios2_p3_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_3_s1_readdata,        --                    .readdata
			out_port   => hex_3_export                                -- external_connection.export
		);

	hex_4 : component nios2_p3_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_4_s1_readdata,        --                    .readdata
			out_port   => hex_4_export                                -- external_connection.export
		);

	hex_5 : component nios2_p3_hex_0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hex_5_s1_address,           --                  s1.address
			write_n    => mm_interconnect_0_hex_5_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_0_hex_5_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_0_hex_5_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_0_hex_5_s1_readdata,          --                    .readdata
			out_port   => hex_5_export                                  -- external_connection.export
		);

	onchip_mem : component nios2_p3_onchip_mem
		port map (
			clk        => clk_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	switch : component nios2_p3_switch
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_switch_s1_readdata,     --                    .readdata
			in_port  => switch_export                             -- external_connection.export
		);

	sysid : component nios2_p3_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component nios2_p3_mm_interconnect_0
		port map (
			clk_clk_clk                             => clk_clk,                                           --                           clk_clk.clk
			cpu_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                    --   cpu_reset_reset_bridge_in_reset.reset
			hex_5_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                -- hex_5_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                 => cpu_data_master_address,                           --                   cpu_data_master.address
			cpu_data_master_waitrequest             => cpu_data_master_waitrequest,                       --                                  .waitrequest
			cpu_data_master_byteenable              => cpu_data_master_byteenable,                        --                                  .byteenable
			cpu_data_master_read                    => cpu_data_master_read,                              --                                  .read
			cpu_data_master_readdata                => cpu_data_master_readdata,                          --                                  .readdata
			cpu_data_master_write                   => cpu_data_master_write,                             --                                  .write
			cpu_data_master_writedata               => cpu_data_master_writedata,                         --                                  .writedata
			cpu_data_master_debugaccess             => cpu_data_master_debugaccess,                       --                                  .debugaccess
			cpu_instruction_master_address          => cpu_instruction_master_address,                    --            cpu_instruction_master.address
			cpu_instruction_master_waitrequest      => cpu_instruction_master_waitrequest,                --                                  .waitrequest
			cpu_instruction_master_read             => cpu_instruction_master_read,                       --                                  .read
			cpu_instruction_master_readdata         => cpu_instruction_master_readdata,                   --                                  .readdata
			cpu_debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --               cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                                  .write
			cpu_debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                                  .read
			cpu_debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                                  .readdata
			cpu_debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                                  .writedata
			cpu_debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                                  .byteenable
			cpu_debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                                  .waitrequest
			cpu_debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                                  .debugaccess
			hex_0_s1_address                        => mm_interconnect_0_hex_0_s1_address,                --                          hex_0_s1.address
			hex_0_s1_write                          => mm_interconnect_0_hex_0_s1_write,                  --                                  .write
			hex_0_s1_readdata                       => mm_interconnect_0_hex_0_s1_readdata,               --                                  .readdata
			hex_0_s1_writedata                      => mm_interconnect_0_hex_0_s1_writedata,              --                                  .writedata
			hex_0_s1_chipselect                     => mm_interconnect_0_hex_0_s1_chipselect,             --                                  .chipselect
			hex_1_s1_address                        => mm_interconnect_0_hex_1_s1_address,                --                          hex_1_s1.address
			hex_1_s1_write                          => mm_interconnect_0_hex_1_s1_write,                  --                                  .write
			hex_1_s1_readdata                       => mm_interconnect_0_hex_1_s1_readdata,               --                                  .readdata
			hex_1_s1_writedata                      => mm_interconnect_0_hex_1_s1_writedata,              --                                  .writedata
			hex_1_s1_chipselect                     => mm_interconnect_0_hex_1_s1_chipselect,             --                                  .chipselect
			hex_2_s1_address                        => mm_interconnect_0_hex_2_s1_address,                --                          hex_2_s1.address
			hex_2_s1_write                          => mm_interconnect_0_hex_2_s1_write,                  --                                  .write
			hex_2_s1_readdata                       => mm_interconnect_0_hex_2_s1_readdata,               --                                  .readdata
			hex_2_s1_writedata                      => mm_interconnect_0_hex_2_s1_writedata,              --                                  .writedata
			hex_2_s1_chipselect                     => mm_interconnect_0_hex_2_s1_chipselect,             --                                  .chipselect
			hex_3_s1_address                        => mm_interconnect_0_hex_3_s1_address,                --                          hex_3_s1.address
			hex_3_s1_write                          => mm_interconnect_0_hex_3_s1_write,                  --                                  .write
			hex_3_s1_readdata                       => mm_interconnect_0_hex_3_s1_readdata,               --                                  .readdata
			hex_3_s1_writedata                      => mm_interconnect_0_hex_3_s1_writedata,              --                                  .writedata
			hex_3_s1_chipselect                     => mm_interconnect_0_hex_3_s1_chipselect,             --                                  .chipselect
			hex_4_s1_address                        => mm_interconnect_0_hex_4_s1_address,                --                          hex_4_s1.address
			hex_4_s1_write                          => mm_interconnect_0_hex_4_s1_write,                  --                                  .write
			hex_4_s1_readdata                       => mm_interconnect_0_hex_4_s1_readdata,               --                                  .readdata
			hex_4_s1_writedata                      => mm_interconnect_0_hex_4_s1_writedata,              --                                  .writedata
			hex_4_s1_chipselect                     => mm_interconnect_0_hex_4_s1_chipselect,             --                                  .chipselect
			hex_5_s1_address                        => mm_interconnect_0_hex_5_s1_address,                --                          hex_5_s1.address
			hex_5_s1_write                          => mm_interconnect_0_hex_5_s1_write,                  --                                  .write
			hex_5_s1_readdata                       => mm_interconnect_0_hex_5_s1_readdata,               --                                  .readdata
			hex_5_s1_writedata                      => mm_interconnect_0_hex_5_s1_writedata,              --                                  .writedata
			hex_5_s1_chipselect                     => mm_interconnect_0_hex_5_s1_chipselect,             --                                  .chipselect
			onchip_mem_s1_address                   => mm_interconnect_0_onchip_mem_s1_address,           --                     onchip_mem_s1.address
			onchip_mem_s1_write                     => mm_interconnect_0_onchip_mem_s1_write,             --                                  .write
			onchip_mem_s1_readdata                  => mm_interconnect_0_onchip_mem_s1_readdata,          --                                  .readdata
			onchip_mem_s1_writedata                 => mm_interconnect_0_onchip_mem_s1_writedata,         --                                  .writedata
			onchip_mem_s1_byteenable                => mm_interconnect_0_onchip_mem_s1_byteenable,        --                                  .byteenable
			onchip_mem_s1_chipselect                => mm_interconnect_0_onchip_mem_s1_chipselect,        --                                  .chipselect
			onchip_mem_s1_clken                     => mm_interconnect_0_onchip_mem_s1_clken,             --                                  .clken
			switch_s1_address                       => mm_interconnect_0_switch_s1_address,               --                         switch_s1.address
			switch_s1_readdata                      => mm_interconnect_0_switch_s1_readdata,              --                                  .readdata
			sysid_control_slave_address             => mm_interconnect_0_sysid_control_slave_address,     --               sysid_control_slave.address
			sysid_control_slave_readdata            => mm_interconnect_0_sysid_control_slave_readdata     --                                  .readdata
		);

	irq_mapper : component nios2_p3_irq_mapper
		port map (
			clk        => clk_clk,                        --       clk.clk
			reset      => rst_controller_reset_out_reset, -- clk_reset.reset
			sender_irq => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component nios2_p3_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component nios2_p3_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_hex_0_s1_write_ports_inv <= not mm_interconnect_0_hex_0_s1_write;

	mm_interconnect_0_hex_1_s1_write_ports_inv <= not mm_interconnect_0_hex_1_s1_write;

	mm_interconnect_0_hex_2_s1_write_ports_inv <= not mm_interconnect_0_hex_2_s1_write;

	mm_interconnect_0_hex_3_s1_write_ports_inv <= not mm_interconnect_0_hex_3_s1_write;

	mm_interconnect_0_hex_4_s1_write_ports_inv <= not mm_interconnect_0_hex_4_s1_write;

	mm_interconnect_0_hex_5_s1_write_ports_inv <= not mm_interconnect_0_hex_5_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of nios2_p3
